---------------------------------------------------------------------------------------------------
--
-- Title       : No Title
-- Design      : sumador
-- Author      : isaiaschavez.co@gmail.com
-- Company     : utm
--
---------------------------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\sumador\sumador\compile\Pruebafulladder4bits.vhd
-- Generated   : Thu Nov  4 22:38:33 2021
-- From        : c:\My_Designs\sumador\sumador\src\Pruebafulladder4bits.bde
-- By          : Bde2Vhdl ver. 2.6
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;


entity Pruebafulladder4bits is 
end Pruebafulladder4bits;

architecture Pruebafulladder4bits of Pruebafulladder4bits is

begin

end Pruebafulladder4bits;
